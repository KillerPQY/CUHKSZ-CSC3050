`timescale 1ns/1ps

module alu_test;

reg[31:0] i_datain, gr1, gr2;

wire[31:0] c;
wire[2:0] flags;
//wire zero;
//wire overflow;
//wire neg;

alu testalu(i_datain, gr1, gr2, c, flags);

initial
begin

$display("instruction:op:func:  gr1   :  gr2   :   c    : reg_A  : reg_B  : reg_C  : flags  ");
$monitor("   %h:%h: %h :%h:%h:%h:%h:%h:%h:%b",
i_datain, testalu.opcode, testalu.func, gr1, gr2, c, testalu.reg_A, testalu.reg_B, testalu.reg_C, testalu.flags);

//add
#10 i_datain<=32'b000000_00001_00000_00000_00000_100000;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_1001;
$display("add");
$display("instruction:op:func:  gr1   :  gr2   :   c    : reg_A  : reg_B  : reg_C  : flags  ");
#10 i_datain<=32'b000000_00001_00000_00000_00000_100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0001;

// addi
#10 i_datain<=32'b001000_00001_00000_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
$display("addi");
$display("instruction:op:func:  gr1   :  gr2   :   c    : reg_A  : reg_B  : reg_C  : flags  ");
#10 i_datain<=32'b001000_00001_00000_0000000000100010;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0001;

// addu
#10 i_datain<=32'b000000_00001_00000_00000_00000_100001;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_1001;
$display("addu");
$display("instruction:op:func:  gr1   :  gr2   :   c    : reg_A  : reg_B  : reg_C  : flags  ");
#10 i_datain<=32'b000000_00001_00000_00000_00000_100001;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0001;

// addiu
#10 i_datain<=32'b001001_00001_00000_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
$display("addiu");
$display("instruction:op:func:  gr1   :  gr2   :   c    : reg_A  : reg_B  : reg_C  : flags  ");
#10 i_datain<=32'b001001_00001_00000_1000000000100000;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0011;

// sub
#10 i_datain<=32'b000000_00001_00000_00000_00000_100010;
gr1<=32'b1111_0000_0000_0000_0000_0000_0101_1101;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
$display("sub");
$display("instruction:op:func:  gr1   :  gr2   :   c    : reg_A  : reg_B  : reg_C  : flags  ");
#10 i_datain<=32'b000000_00001_00000_00000_00000_100010;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b0111_0000_0000_0000_0000_0000_0101_1101;

// subu
#10 i_datain<=32'b000000_00001_00000_00000_00000_100011;
gr1<=32'b0111_0000_0000_0000_0000_0000_0101_1101;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
$display("subu");
$display("instruction:op:func:  gr1   :  gr2   :   c    : reg_A  : reg_B  : reg_C  : flags  ");
#10 i_datain<=32'b000000_00001_00000_00000_00000_100011;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b0111_0000_0000_0000_0000_0000_0101_1101;

// and
#10 i_datain<=32'b000000_00001_00000_00000_00000_100100;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;
$display("and");
$display("instruction:op:func:  gr1   :  gr2   :   c    : reg_A  : reg_B  : reg_C  : flags  ");
#10 i_datain<=32'b000000_00001_00000_00000_00000_100100;
gr1<=32'b1000_0000_1001_0000_0000_0000_0000_0000;
gr2<=32'b0000_0000_1001_0000_0000_0000_0011_0010;

// andi
#10 i_datain<=32'b001100_00001_00000_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
$display("andi");
$display("instruction:op:func:  gr1   :  gr2   :   c    : reg_A  : reg_B  : reg_C  : flags  ");
#10 i_datain<=32'b001100_00001_00000_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0010_0000;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0001;

// nor
#10 i_datain<=32'b000000_00001_00000_00000_00000_100111;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;
$display("nor");
$display("instruction:op:func:  gr1   :  gr2   :   c    : reg_A  : reg_B  : reg_C  : flags  ");
#10 i_datain<=32'b000000_00001_00000_00000_00000_100111;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0011_0010;

// or
#10 i_datain<=32'b000000_00001_00000_00000_00000_100101;
gr1<=32'b1111_1100_0010_0000_0000_0000_0000_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0011_0010;
$display("or");
$display("instruction:op:func:  gr1   :  gr2   :   c    : reg_A  : reg_B  : reg_C  : flags  ");
#10 i_datain<=32'b000000_00001_00000_00000_00000_100101;
gr1<=32'b0100_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;

// ori
#10 i_datain<=32'b001101_00001_00000_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
$display("ori");
$display("instruction:op:func:  gr1   :  gr2   :   c    : reg_A  : reg_B  : reg_C  : flags  ");
#10 i_datain<=32'b001101_00001_00000_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0010_0000;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0001;

// xor
#10 i_datain<=32'b000000_00001_00000_00000_00000_100110;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;
$display("xor");
$display("instruction:op:func:  gr1   :  gr2   :   c    : reg_A  : reg_B  : reg_C  : flags  ");
#10 i_datain<=32'b000000_00001_00000_00000_00000_100110;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0011_0010;

// xori
#10 i_datain<=32'b001110_00001_00000_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
$display("xori");
$display("instruction:op:func:  gr1   :  gr2   :   c    : reg_A  : reg_B  : reg_C  : flags  ");
#10 i_datain<=32'b001110_00001_00000_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0010_0000;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0001;

// beq
#10 i_datain<=32'b000100_00001_00000_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
$display("beq");
$display("instruction:op:func:  gr1   :  gr2   :   c    : reg_A  : reg_B  : reg_C  : flags  ");
#10 i_datain<=32'b000100_00001_00000_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0010_0000;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0001;

// bne
#10 i_datain<=32'b000101_00001_00000_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
$display("bne");
$display("instruction:op:func:  gr1   :  gr2   :   c    : reg_A  : reg_B  : reg_C  : flags  ");
#10 i_datain<=32'b000101_00001_00000_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0010_0000;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0001;

// slt
#10 i_datain<=32'b000000_00001_00000_00000_00000_101010;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;
$display("slt");
$display("instruction:op:func:  gr1   :  gr2   :   c    : reg_A  : reg_B  : reg_C  : flags  ");
#10 i_datain<=32'b000000_00001_00000_00000_00000_101010;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0011_0010;

// slti
#10 i_datain<=32'b001010_00001_00000_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
$display("slti");
$display("instruction:op:func:  gr1   :  gr2   :   c    : reg_A  : reg_B  : reg_C  : flags  ");
#10 i_datain<=32'b001010_00001_00000_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0010_0000;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0001;

// sltiu
#10 i_datain<=32'b001011_00001_00000_0000000000100000;
gr1<=32'b0000_0000_0000_0000_0000_0000_0010_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
$display("stliu");
$display("instruction:op:func:  gr1   :  gr2   :   c    : reg_A  : reg_B  : reg_C  : flags  ");
#10 i_datain<=32'b001011_00001_00000_0000000000010000;
gr1<=32'b0000_0000_0000_0000_0000_0000_0010_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0001;

// sltu
#10 i_datain<=32'b000000_00001_00000_00000_00000_101011;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;
$display("sltu");
$display("instruction:op:func:  gr1   :  gr2   :   c    : reg_A  : reg_B  : reg_C  : flags  ");
#10 i_datain<=32'b000000_00001_00000_00000_00000_101011;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0011_0010;

// lw
#10 i_datain<=32'b100011_00001_00000_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
$display("lw");
$display("instruction:op:func:  gr1   :  gr2   :   c    : reg_A  : reg_B  : reg_C  : flags  ");
#10 i_datain<=32'b100011_00001_00000_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0010_0000;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0001;

// sw
#10 i_datain<=32'b101011_00001_00000_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
$display("sw");
$display("instruction:op:func:  gr1   :  gr2   :   c    : reg_A  : reg_B  : reg_C  : flags  ");
#10 i_datain<=32'b101011_00001_00000_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0010_0000;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0001;

// sll
#10 i_datain<=32'b000000_00001_00000_00000_00001_000000;
gr1<=32'b1111_1100_0010_0000_0000_0000_0000_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
$display("sll");
$display("instruction:op:func:  gr1   :  gr2   :   c    : reg_A  : reg_B  : reg_C  : flags  ");
#10 i_datain<=32'b000000_00001_00000_00000_00000_000000;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0100;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;

// sllv
#10 i_datain<=32'b000000_00001_00000_00000_00000_000100;
gr1<=32'b0000_0000_0000_0000_0000_0000_0010_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0011_0010;
$display("sllv");
$display("instruction:op:func:  gr1   :  gr2   :   c    : reg_A  : reg_B  : reg_C  : flags  ");
#10 i_datain<=32'b000000_00001_00000_00000_00000_000100;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0110;
gr2<=32'b0000_0000_0000_0000_0000_0000_0001_0000;

// srl
#10 i_datain<=32'b000000_00001_00000_00000_00001_000010;
gr1<=32'b1111_1100_0010_0000_0000_0000_0000_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
$display("srl");
$display("instruction:op:func:  gr1   :  gr2   :   c    : reg_A  : reg_B  : reg_C  : flags  ");
#10 i_datain<=32'b000000_00001_00000_00000_00000_000010;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0100;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;

// srlv
#10 i_datain<=32'b000000_00001_00000_00000_00000_000110;
gr1<=32'b0000_0000_0000_0000_0000_0000_0010_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0011_0010;
$display("srlv");
$display("instruction:op:func:  gr1   :  gr2   :   c    : reg_A  : reg_B  : reg_C  : flags  ");
#10 i_datain<=32'b000000_00001_00000_00000_00000_000110;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0110;
gr2<=32'b0000_0000_0000_0000_0000_0000_0001_0000;

// sra
#10 i_datain<=32'b000000_00001_00000_00000_00001_000011;
gr1<=32'b1111_1100_0010_0000_0000_0000_0000_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0011_0010;
$display("sra");
$display("instruction:op:func:  gr1   :  gr2   :   c    : reg_A  : reg_B  : reg_C  : flags  ");
#10 i_datain<=32'b000000_00001_00000_00000_00001_000011;
gr1<=32'b0100_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;

// srav
#10 i_datain<=32'b000000_00001_00000_00000_00000_000110;
gr1<=32'b0000_0000_0000_0000_0000_0000_0010_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0011_0010;
$display("srav");
$display("instruction:op:func:  gr1   :  gr2   :   c    : reg_A  : reg_B  : reg_C  : flags  ");
#10 i_datain<=32'b000000_00001_00000_00000_00000_000110;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0110;
gr2<=32'b0000_0000_0000_0000_0000_0000_0001_0000;


#10 $finish;
end
endmodule