`include "CPU.v"

`timescale 100fs/100fs

module test_CPU;
CPU CPU_1();
endmodule